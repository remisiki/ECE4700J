module arbiterFSM(
        input clock, reset, A, B,
        output grant_to_A, grant_to_B
        ); 

//TODO: Start your design here

endmodule